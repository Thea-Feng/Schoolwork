`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain, gr1, gr2;


wire[31:0] c;
wire[2:0] flags;

alu test(i_datain,gr1, gr2, c, flags);

initial
begin

$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
$monitor("   %h:%h: %h :%h:%h:%h:%h:%h:   %h  :     %h    :     %h",
i_datain, test.opcode, test.func, gr1 , gr2, test.reg_A, test.reg_B, test.c, test.zero, test.neg, test.overflow);

//add
#10 i_datain<=32'b000000_00000_00001_00010_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b0000_0000_0000_0000_0000_0000_0001_0001;
$display("add");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_1001;
gr2<=32'b1000_0000_0000_0000_0000_0000_1000_0110;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100000;
gr1<=32'b0100_0000_0000_0000_0000_0000_0110_0010;
gr2<=32'b0100_0000_0000_0000_0000_0000_0011_0001;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_1101_1101;
gr2<=32'b1111_1111_1111_1111_1111_1111_0010_0011;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0101_1101;
gr2<=32'b1111_1111_1111_1111_1111_1111_0010_0011;

//addi
#10 i_datain<=32'b001000_00000_00001_1000000000100011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("addi");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001000_00000_00001_0000000100100010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;

#10 i_datain<=32'b001000_00000_00001_0000111000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;

#10 i_datain<=32'b001000_00000_00001_1110000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0001;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

//addu
#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
$display("addu");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0100_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b0000_0000_0000_0000_0000_0000_1101_1101;
gr2<=32'b1111_1111_1111_1111_1111_1111_0010_0011;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0101_1101;
gr2<=32'b1111_1111_1111_1111_1111_1111_0010_0011;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//addiu
#10 i_datain<=32'b001001_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("addiu");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001001_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

#10 i_datain<=32'b001001_00000_00001_0000000000000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//sub
#10 i_datain<=32'b000000_00000_00001_00010_00000_100010;
gr1<=32'b1111_0000_0000_0000_0000_0000_0101_1101;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("sub");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b0111_0000_0000_0000_0000_0000_0101_1101;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100010;
gr1<=32'b0000_0000_0000_0000_0010_0000_0000_0001;
gr2<=32'b1111_0000_0000_1101_0000_0000_0101_1101;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100010;
gr1<=32'b0000_1111_0000_0000_0000_1111_0000_0000;
gr2<=32'b0000_1111_0000_0000_0000_1111_0000_0000;

//subu
#10 i_datain<=32'b000000_00000_00001_00010_00000_100011;
gr1<=32'b0111_0000_0000_0000_1110_0000_0101_1101;
gr2<=32'b1000_0000_1111_0000_0000_0000_0000_0001;
$display("subu");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0111_0000_0000_0000_0000_0000_0101_1101;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100011;
gr1<=32'b0000_0001_0000_0111_0000_0000_0000_0001;
gr2<=32'b1111_0011_0000_0000_1110_0000_0101_1101;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100011;
gr1<=32'b0000_0000_0000_0000_1100_1000_0000_0001;
gr2<=32'b0000_0000_0011_0000_0000_0011_0101_1101;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100011;
gr1<=32'b0000_0000_0000_0000_0000_0011_0000_0000;
gr2<=32'b0000_0000_1100_0000_0000_0000_0000_0000;

//and
#10 i_datain<=32'b000000_00000_00001_00010_00000_100100;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("and");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100100;
gr1<=32'b1000_0000_1001_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_1001_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100100;
gr1<=32'b1000_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100100;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//andi
#10 i_datain<=32'b001100_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("andi");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001100_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b001100_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//nor
#10 i_datain<=32'b000000_00000_00001_00010_00000_100111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("nor");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100111;
gr1<=32'b1000_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//or
#10 i_datain<=32'b000000_00000_00001_00010_11000_100101;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;
$display("or");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_100101;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

#10 i_datain<=32'b000000_00000_00001_00010_11000_100101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//ori
#10 i_datain<=32'b001101_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("ori");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001101_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b001101_00000_00001_0000000000000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//xor
#10 i_datain<=32'b000000_00000_00001_00010_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("xor");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100110;
gr1<=32'b1000_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//xori
#10 i_datain<=32'b001110_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("xori");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001110_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b001110_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//beq/bne
#10 i_datain<=32'b000100_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("beq/bne");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000100_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b000100_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//slt
#10 i_datain<=32'b000000_00000_00001_00010_00000_101010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("slt");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_101010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_101010;
gr1<=32'b0100_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_101010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//slti
#10 i_datain<=32'b001010_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("slti");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001010_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b001010_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//sltu
#10 i_datain<=32'b000000_00000_00001_00010_00000_101011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
$display("sltu");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_00000_101011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_101011;
gr1<=32'b1000_1100_0010_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b000000_00000_00001_00010_00000_101011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//stliu
#10 i_datain<=32'b001011_00000_00001_0000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
$display("stliu");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b001011_00000_00001_0000000000010000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b001011_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;

#10 i_datain<=32'b001011_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//sw
#10 i_datain<=32'b101011_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0111;
$display("sw");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b101011_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0001;

#10 i_datain<=32'b101011_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//lw
#10 i_datain<=32'b100011_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0010_0000_0111;
gr2<=32'b1000_0000_0000_0000_0000_0010_0000_0111;
$display("lw");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b100011_00000_00001_1000000000100000;
gr1<=32'b1000_0000_0000_0000_0000_0011_0010_0000;
gr2<=32'b1000_0000_0000_0000_0011_0000_0000_0001;

#10 i_datain<=32'b100011_00000_00001_1000000000100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0011_0001;
gr2<=32'b0000_0000_0000_0000_0011_0000_0000_0011;

//sll
#10 i_datain<=32'b000000_00000_00001_00010_11000_000000;
gr1<=32'b1111_1100_0010_0000_0011_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0011_0011_0010;
$display("sll");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//sllv
#10 i_datain<=32'b000000_00000_00001_00010_11000_000100;
gr2<=32'b0000_0000_0000_0000_0000_0011_0010_0000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
$display("sllv");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000100;
gr2<=32'b0000_0000_0000_0011_0000_0000_0000_0110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//srl
#10 i_datain<=32'b000000_00000_00001_00010_11000_000010;
gr1<=32'b1111_1100_0010_0100_0000_0000_0000_0000;
gr2<=32'b0000_0000_0100_0000_0000_0010_0011_0010;
$display("srl");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000010;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//srlv
#10 i_datain<=32'b000000_00000_00001_00010_11000_000110;
gr2<=32'b0000_0000_0000_0000_0010_0000_0010_0000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
$display("srlv");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000110;
gr2<=32'b1000_0000_0000_0100_0010_0000_0000_0110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1001;

//sra
#10 i_datain<=32'b000000_00000_00001_00010_11000_000011;
gr1<=32'b1111_1100_0010_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0011;
$display("sra");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000011;
gr1<=32'b0100_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//srav
#10 i_datain<=32'b000000_00000_00001_00010_11000_000111;
gr2<=32'b1000_0000_0100_0000_0010_0000_0010_0001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0001_0011;
$display("srav");
$display("instruction:op:func:  gr1   :  gr2   : reg_A  : reg_B  : reg_C  : zero : negative : overflow");
#10 i_datain<=32'b000000_00000_00001_00010_11000_000111;
gr2<=32'b0000_0000_0000_0010_0001_0000_0000_0111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0001_0010;

//invalid input
#10 i_datain<=32'b111111_00000_00001_00010_11000_000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0010_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0011_0010;

#10 i_datain<=32'b101111_00000_00001_00010_11000_000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0110;
gr2<=32'b1111_1111_1101_1111_1111_1111_1111_1101;






#10 $finish;
end
endmodule
